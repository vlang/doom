[translated]
module main

[typedef]
struct C.FILE {}

// vstart

const ( // empty enum
)

[c: 'A_Light0']
fn a_light0()

[c: 'A_WeaponReady']
fn a_weaponready()

[c: 'A_Lower']
fn a_lower()

[c: 'A_Raise']
fn a_raise()

[c: 'A_Punch']
fn a_punch()

[c: 'A_ReFire']
fn a_refire()

[c: 'A_FirePistol']
fn a_firepistol()

[c: 'A_Light1']
fn a_light1()

[c: 'A_FireShotgun']
fn a_fireshotgun()

[c: 'A_Light2']
fn a_light2()

[c: 'A_FireShotgun2']
fn a_fireshotgun2()

[c: 'A_CheckReload']
fn a_checkreload()

[c: 'A_OpenShotgun2']
fn a_openshotgun2()

[c: 'A_LoadShotgun2']
fn a_loadshotgun2()

[c: 'A_CloseShotgun2']
fn a_closeshotgun2()

[c: 'A_FireCGun']
fn a_firecgun()

[c: 'A_GunFlash']
fn a_gunflash()

[c: 'A_FireMissile']
fn a_firemissile()

[c: 'A_Saw']
fn a_saw()

[c: 'A_FirePlasma']
fn a_fireplasma()

[c: 'A_BFGsound']
fn a_bfgsound()

[c: 'A_FireBFG']
fn a_firebfg()

[c: 'A_BFGSpray']
fn a_bfgspray()

[c: 'A_Explode']
fn a_explode()

[c: 'A_Pain']
fn a_pain()

[c: 'A_PlayerScream']
fn a_playerscream()

[c: 'A_Fall']
fn a_fall()

[c: 'A_XScream']
fn a_xscream()

[c: 'A_Look']
fn a_look()

[c: 'A_Chase']
fn a_chase()

[c: 'A_FaceTarget']
fn a_facetarget()

[c: 'A_PosAttack']
fn a_posattack()

[c: 'A_Scream']
fn a_scream()

[c: 'A_SPosAttack']
fn a_sposattack()

[c: 'A_VileChase']
fn a_vilechase()

[c: 'A_VileStart']
fn a_vilestart()

[c: 'A_VileTarget']
fn a_viletarget()

[c: 'A_VileAttack']
fn a_vileattack()

[c: 'A_StartFire']
fn a_startfire()

[c: 'A_Fire']
fn a_fire()

[c: 'A_FireCrackle']
fn a_firecrackle()

[c: 'A_Tracer']
fn a_tracer()

[c: 'A_SkelWhoosh']
fn a_skelwhoosh()

[c: 'A_SkelFist']
fn a_skelfist()

[c: 'A_SkelMissile']
fn a_skelmissile()

[c: 'A_FatRaise']
fn a_fatraise()

[c: 'A_FatAttack1']
fn a_fatattack1()

[c: 'A_FatAttack2']
fn a_fatattack2()

[c: 'A_FatAttack3']
fn a_fatattack3()

[c: 'A_BossDeath']
fn a_bossdeath()

[c: 'A_CPosAttack']
fn a_cposattack()

[c: 'A_CPosRefire']
fn a_cposrefire()

[c: 'A_TroopAttack']
fn a_troopattack()

[c: 'A_SargAttack']
fn a_sargattack()

[c: 'A_HeadAttack']
fn a_headattack()

[c: 'A_BruisAttack']
fn a_bruisattack()

[c: 'A_SkullAttack']
fn a_skullattack()

[c: 'A_Metal']
fn a_metal()

[c: 'A_SpidRefire']
fn a_spidrefire()

[c: 'A_BabyMetal']
fn a_babymetal()

[c: 'A_BspiAttack']
fn a_bspiattack()

[c: 'A_Hoof']
fn a_hoof()

[c: 'A_CyberAttack']
fn a_cyberattack()

[c: 'A_PainAttack']
fn a_painattack()

[c: 'A_PainDie']
fn a_paindie()

[c: 'A_KeenDie']
fn a_keendie()

[c: 'A_BrainPain']
fn a_brainpain()

[c: 'A_BrainScream']
fn a_brainscream()

[c: 'A_BrainDie']
fn a_braindie()

[c: 'A_BrainAwake']
fn a_brainawake()

[c: 'A_BrainSpit']
fn a_brainspit()

[c: 'A_SpawnSound']
fn a_spawnsound()

[c: 'A_SpawnFly']
fn a_spawnfly()

[c: 'A_BrainExplode']
fn a_brainexplode()
