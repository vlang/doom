[translated]
module main

[typedef]
struct C.FILE {}

// vstart
