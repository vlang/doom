[translated]
module main


[typedef]
struct C.FILE {}


// vstart


const ( // empty enum
)

// skipped extern global gamevariant
[weak]__global ( gamedescription &i8 

)

[weak]__global ( modifiedgame bool 

)

/*!*/[weak] __global ( gamevariant  = GameVariant_t (GameVariant_t.vanilla)
)

